// Entry point for examples using imgui.
// Import the example you want and call its main

module main

// Note, flags are loaded on import
import examples.glfw_vulkan


fn main() {
  glfw_vulkan.main()
}
